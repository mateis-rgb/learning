* AC Analysis, 1k lowPass, 4th order Butterworth, 2 stages using AD711

* Input signal for AC and transient sinusoidal analysis
VIN IN 0 AC 1 DC 0 SINE(0 1.06 100)
* VNOISE IN 0 AC 0 DC 0

XA IN OUTA VCCG VEEG 0 sallenKeylowPassStageA
XB OUTA OUT VCCG VEEG 0 sallenKeylowPassStageB

VP VCCG 0 5
VM VEEG 0 -5

*Simulation directive lines for AC Analysis
.AC DEC 100 100 20k
*.TRAN 1n 3.99m
*.NOISE V(OUT) VNOISE DEC 100 100 20k
.PROBE

.SUBCKT sallenKeylowPassStageA IN OUT VCC VEE GND
X1 INP OUT VCC VEE OUT AD711
R1 IN 1 26.7k
R2 1 INP 95.3k
C1 1 OUT 10n
C2 INP GND 1n
.ENDS sallenKeylowPassStageA

.SUBCKT sallenKeylowPassStageB IN OUT VCC VEE GND
X1 INP OUT VCC VEE OUT AD711
R1 IN 1 100k
R2 1 INP 191k
C1 1 OUT 1.3n
C2 INP GND 1n
.ENDS sallenKeylowPassStageB

* AD711 SPICE Macro-model  
* Description: Amplifier 
* Generic Desc: 10/30V, BIP, OP, Fast, Precision, 1X
* Developed by: JLW / PMI, TRW / ADI
* Revision History: 08/10/2012 - Updated to new header style
* 3.0 (03/1991) - Corrected VOS to be 0.1mV.
* Copyright 1991, 2012 by Analog Devices.
*
* Refer to http://www.analog.com/Analog_Root/static/techSupport/designTools/spiceModels/license/spice_general.html for License Statement. Use of this model
* indicates your acceptance with the terms and provisions in the License Statement.
*
* BEGIN Notes:
*
* Not Modeled:
*
* Parameters modeled include:
* This version of the AD711 model simulates the typical 
* parameters corresponding to the device data sheet.
*
* END Notes
*
* Node assignments
* connections: non-inverting input 
*              |  inverting input  
*              |  |  positive supply
*              |  |  |  negative supply
*              |  |  |  |  output
*              |  |  |  |  |
.SUBCKT AD711 13 15 12 16 14
* 
VOS 15 8 DC 0.1E-3
EC 9 0 (14,0) 1
C1 6 7 .5E-12
RP 16 12 12E3
GB 11 0 (3,0) 1.67E3
RD1 6 16 16E3
RD2 7 16 16E3
ISS 12 1 DC 100E-6
CCI 3 11 150E-12
GCM 0 3 (0,1) 1.76E-9
GA 3 0 (7,6) 2.3E-3
RE 1 0 2.5E6
RGM 3 0 1.69E3
VC 12 2 DC 2.8
VE 10 16 DC 2.8
RO1 11 14 25
CE 1 0 2E-12
RO2 0 11 30
RS1 1 4 5.77E3
RS2 1 5 5.77E3
J1 6 13 4 FET
J2 7 8 5 FET
DC 14 2 DIODE
DE 10 14 DIODE
DP 16 12 DIODE
D1 9 11 DIODE
D2 11 9 DIODE
IOS 15 13 5E-12
.MODEL DIODE D()
.MODEL FET PJF(VTO=-1 BETA=1E-3 IS=15E-12)
.ENDS


